module k14(output [48:1] out);
    assign out = 48'b110100111010100010101100100110000000000110101100;
endmodule
