module k2(output [48:1] out);
    assign out = 48'b001000001011111010100010101000001100000000010111;
endmodule
